library UNISIM;
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use UNISIM.VComponents.all;

entity N1 is
end N1;

architecture Behavioral of N1 is

begin


end Behavioral;

