library ieee;use ieee.std_logic_1164.all;entity tff is	port (Rst, clk, T : in ustd_logic := '1';		     Q : out std_ulogic);end tff;architecture behave of tff isbegin	process (Rst, clk) is	variable qtmp :std_ulogic;	begin		if (Rst = '1') then		   qtmp := '0';		elsif rising_edge( clk) then		    if T = '1' then		       qtmp := not qtmp;		    end if;	       end if;	Q <= qtmp;	end process;end behave; 	